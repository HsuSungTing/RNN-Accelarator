`timescale 1ns / 0.1ps
module test_exam;
    reg [31:0]FP_A,FP_B;
    wire [31:0]FP_out;

    MUT U1(.FP_A(FP_A),.FP_B(FP_B),.FP_out(FP_out));

    initial begin
        FP_A=32'b01000000001001110000101000111101;//2.61，確定是2.61
        FP_B=32'b00111110100101000111101011100001;//0.29，確定是0.29
        
        #5
        FP_A=32'b00111111110001111010111000010100;//1.56。確定是1.56
        FP_B=32'b00111111100111010111000010100100;//1.23，確定是1.23

        #5
        FP_A=32'b01000011000000111000111101011100;//131.56。確定
        FP_B=32'b01000011011010101100011110101110;//234.78，確定

        #5
        FP_A=32'b00111111110001111010111000010100;//131.56。確定
        FP_B=32'b00111111101011110101110000101001;//234.78，確定
        
    end

endmodule