`timescale 1ns / 0.1ps
module test_exam;
    reg  [31:0]FP_A,FP_B;
    wire [31:0]FP_out;

    ADD U0(.FP_A(FP_A),.FP_B(FP_B),.FP_out(FP_out));

    initial begin
        FP_A=32'b01000101010010111000010100011111;    //3256.32
        FP_B=32'b00111110011101011100001010001111;    //0.24
        
        #5
        FP_A=32'b10111111101010001111010111000011;    //-1.32
        FP_B=32'b11000000001000101000111101011100;    //-2.54
        //answer=11000000011101110000101000111101

        #5
        FP_A=32'b0011_1111_0100_0001_1100_0100_0011_0001;    //-1.32
        FP_B=32'b0011_1111_1111_0101_1001_1011_0011_1100;    //-2.54
        //answer=11000000011101110000101000111101
    end

endmodule