`timescale 1ns / 0.1ps
module test_exam;
    reg  clk, rst_n, in_valid;
    reg [31:0] weight_u, weight_w, weight_v, data_x, data_h;
    wire out_valid;

    RNN T0(.clk(clk),.rst_n(rst_n),.in_valid(in_valid),.weight_u(weight_u),.weight_w(weight_w),.weight_v(weight_v),
    .data_x(data_x),.data_h(data_h),.out_valid(out_valid),.out(out));

    always 
        #5 clk=~clk;
    initial begin
        rst_n=1'b0;clk=1'b0;in_valid=1'b0;
        #5 rst_n=1'b1;in_valid=1'b0;
        #5 rst_n=1'b0;in_valid=1'b0;
        #5 in_valid=1'b0;
        #10 in_valid=1'b1;weight_u=32'b01000000001001110000101000111101;weight_w=32'b00111111000011110101110000101001;weight_v=32'b01000000001000000000000000000000;data_x=32'b00111110100101000111101011100001;data_h=32'b00111111100111000010100011110110;
        #10 weight_u=32'b00111111110001111010111000010100;weight_w=32'b01000000000100010100011110101110;weight_v=32'b00111111001000010100011110101110;data_x=32'b00111111100111010111000010100100;data_h=32'b00111110000001010001111010111000;
        #10 weight_u=32'b01000000000100010100011110101110;weight_w=32'b00111111001111010111000010100100;weight_v=32'b00111111010001010001111010111000;data_x=32'b00111111101011110101110000101001;data_h=32'b01000000001000111101011100001010;

        #10 weight_u=32'b00111111010100011110101110000101;weight_w=32'b00111111111001100110011001100110;weight_v=32'b00111111011110000101000111101100;data_x=32'b00111101101000111101011100001010;
        #10 weight_u=32'b01000000000101110000101000111101;weight_w=32'b00111111000010100011110101110001;weight_v=32'b00111111001010001111010111000011;data_x=32'b00111111100011001100110011001101;
        #10 weight_u=32'b00111110001011100001010001111011;weight_w=32'b01000000000000011110101110000101;weight_v=32'b01000000001101011100001010001111;data_x=32'b00111111101101110000101000111101;

        #10 weight_u=32'b01000000001010000101000111101100;weight_w=32'b01000000000110101110000101001000;weight_v=32'b01000000000111010111000010100100;data_x=32'b00111111110100011110101110000101;
        #10 weight_u=32'b01000000000010100011110101110001;weight_w=32'b00111110010011001100110011001101;weight_v=32'b00111111111101000111101011100001;data_x=32'b01000000001110101110000101001000;
        #10 weight_u=32'b00111111110001111010111000010100;weight_w=32'b00111111011110000101000111101100;weight_v=32'b00111111010000101000111101011100;data_x=32'b01000000000011110101110000101001;
       
    end

endmodule