`timescale 1ns / 0.1ps
module test_exam;
    reg [31:0]M_00,M_01,M_02,M_10,M_11,M_12,M_20,M_21,M_22;
    reg [31:0]in_0,in_1,in_2;

    wire [31:0]Sum_row0,Sum_row1,Sum_row2;

    matrix_MUT U0(.M_00(M_00),.M_01(M_01),.M_02(M_02),
    .M_10(M_10),.M_11(M_11),.M_12(M_12),
    .M_20(M_20),.M_21(M_21),.M_22(M_22),
    .in_0(in_0),.in_1(in_1),.in_2(in_2),
    .Sum_row0(Sum_row0),.Sum_row1(Sum_row1),.Sum_row2(Sum_row2));

    initial begin
        M_00=32'b01000000001001110000101000111101;//2.61
        M_01=32'b00111111110001111010111000010100;//1.56
        M_02=32'b01000000000100010100011110101110;//2.27
        M_10=32'b00111111010100011110101110000101;//0.82
        M_11=32'b01000000000101110000101000111101;//2.36
        M_12=32'b00111110001011100001010001111011;//0.17
        M_20=32'b01000000001010000101000111101100;//2.63
        M_21=32'b01000000000010100011110101110001;//2.16
        M_22=32'b00111111110001111010111000010100;//1.56
        
        in_0=32'b00111110100101000111101011100001;//0.29
        in_1=32'b00111111100111010111000010100100;//1.23
        in_2=32'b00111111101011110101110000101001;//1.37
        
    end
endmodule
